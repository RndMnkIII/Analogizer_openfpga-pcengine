// unnamed.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module unnamed (
		input  wire  inclk1x,   //  altclkctrl_input.inclk1x
		input  wire  inclk0x,   //                  .inclk0x
		input  wire  clkselect, //                  .clkselect
		output wire  outclk     // altclkctrl_output.outclk
	);

	unnamed_altclkctrl_0 altclkctrl_0 (
		.inclk1x   (inclk1x),   //  altclkctrl_input.inclk1x
		.inclk0x   (inclk0x),   //                  .inclk0x
		.clkselect (clkselect), //                  .clkselect
		.outclk    (outclk)     // altclkctrl_output.outclk
	);

endmodule
